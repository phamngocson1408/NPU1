`timescale 100ps / 1ps
`define CYCLE 		20
`define RUN_TIME	10


`define CHANNEL_STACKING

`ifdef CHANNEL_STACKING
	`undef CHANNEL_PADDING
`else
	`define CHANNEL_PADDING
`endif

//`define COMB_DAT_CHUNK

`ifdef CHANNEL_STACKING
	`define COMB_DAT_CHUNK
`endif

`ifdef CHANNEL_STACKING
	`define CHUNK_SIZE	128*2	//Bytes
`elsif CHANNEL_PADDING
	`define CHUNK_SIZE	128	//Bytes
`endif

`define BUS_SIZE		8	//Bytes
`define PREFIX_SUM_SIZE		8	//bits
`define OUTPUT_BUF_SIZE		32	//bits
`define COMPUTE_UNIT_NUM	1
`define DAT_SIZE		8	//bits 
`define DIVIDED_CHANNEL_NUM 	8

`define IFM_DENSE_RATE 		70
`define FILTER_DENSE_RATE 	70

// Do not change when FULL_CHANNEL and CHANNEL_PADDING
`define LAYER_CHANNEL_NUM_MAX 	192
`define LAYER_FILTER_SIZE_MAX 	5
`define LAYER_OUTPUT_SIZE_MAX 	10
`define LAYER_IFM_SIZE_MAX 	(`LAYER_FILTER_SIZE_MAX + `LAYER_OUTPUT_SIZE_MAX - 1)

`define LAYER_CHANNEL_NUM 	128
`define LAYER_FILTER_SIZE_X 	4
`define LAYER_FILTER_SIZE_Y 	4
`define LAYER_OUTPUT_SIZE_X 	4
`define LAYER_OUTPUT_SIZE_Y 	4
`define LAYER_IFM_SIZE_X 	(`LAYER_FILTER_SIZE_X + `LAYER_OUTPUT_SIZE_X - 1)
`define LAYER_IFM_SIZE_Y 	(`LAYER_FILTER_SIZE_Y + `LAYER_OUTPUT_SIZE_Y - 1)

`define OUTPUT_BUF_NUM		(`LAYER_OUTPUT_SIZE_Y * `LAYER_OUTPUT_SIZE_X) 

`ifdef CHANNEL_STACKING
	`define SRAM_IFM_NUM 		((`LAYER_CHANNEL_NUM / `DIVIDED_CHANNEL_NUM) * `LAYER_IFM_SIZE_Y)
	`define SRAM_FILTER_NUM 	((`LAYER_CHANNEL_NUM / `DIVIDED_CHANNEL_NUM) * `COMPUTE_UNIT_NUM)
`elsif CHANNEL_PADDING
	`define SRAM_IFM_NUM 		(2 * (`LAYER_IFM_SIZE_Y * `LAYER_IFM_SIZE_X))
	`define SRAM_FILTER_NUM 	(2 * (`LAYER_FILTER_SIZE_Y * `LAYER_FILTER_SIZE_X) * `COMPUTE_UNIT_NUM)
`endif

`define WR_DAT_CYC_NUM		(`CHUNK_SIZE/`BUS_SIZE)
`define RD_DAT_CYC_NUM		(`CHUNK_SIZE/`PREFIX_SUM_SIZE)

`ifdef CHANNEL_STACKING
	`define SIM_CHUNK_SIZE	128*2
`elsif CHANNEL_PADDING
	`define SIM_CHUNK_SIZE	128	//Bytes
`endif

`define SIM_WR_DAT_CYC_NUM	(`SIM_CHUNK_SIZE/`BUS_SIZE)
`define SIM_RD_DAT_CYC_NUM	(`SIM_CHUNK_SIZE/`PREFIX_SUM_SIZE)

//`define SHORT_CHANNEL
//`ifdef SHORT_CHANNEL
//	`undef FULL_CHANNEL
//`else
//	`define FULL_CHANNEL
//`endif


