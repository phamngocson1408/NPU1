`define COMB_DAT_CHUNK