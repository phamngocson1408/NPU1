`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 07/24/2022 06:03:16 PM
// Design Name: 
// Module Name: Data_Chunk
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module Dat_Chunk_Comb #(
	 parameter MEM_SIZE = 128	//Bytes
	,parameter BUS_SIZE = 16	//Bytes
	,parameter PREFIX_SUM_SIZE = 16	//bits	
)(
	 input rst_i
	,input clk_i
	,input [BUS_SIZE-1:0] wr_sparsemap_i
	,input [BUS_SIZE-1:0][7:0] wr_nonzero_data_i 	//Bandwidth = 128 Bytes
	,input wr_valid_i
	,input [$clog2(MEM_SIZE/BUS_SIZE)-1:0] wr_count_i

	,output [MEM_SIZE:1][7:0] rd_nonzero_data_o
	,output logic [MEM_SIZE-1:0] rd_sparsemap_o	
);
	
	logic [MEM_SIZE-1:0] mem_sparsemap_r;
	//The Data array should start from 1
	logic [MEM_SIZE:1][7:0] mem_nonzero_data_r;

	// Write data
	always_ff @(posedge clk_i) begin
		if (rst_i) begin
			mem_sparsemap_r <= #1 {MEM_SIZE{1'b0}};
			mem_nonzero_data_r <= #1 {MEM_SIZE{8'h00}};
		end
		else if (wr_valid_i) begin
			for (integer i=0; i<MEM_SIZE/BUS_SIZE; i=i+1) begin
				if (wr_count_i == i) begin
					mem_sparsemap_r[BUS_SIZE*i +: BUS_SIZE] <= #1 wr_sparsemap_i;
					mem_nonzero_data_r[(BUS_SIZE*i+1) +: BUS_SIZE] <= #1 wr_nonzero_data_i;
				end
			end
		end
	end

	assign rd_nonzero_data_o = mem_nonzero_data_r;
	assign rd_sparsemap_o = mem_sparsemap_r;

endmodule
