//`define COMB_DAT_CHUNK
`define PREFIX_SUM_SIZE 8